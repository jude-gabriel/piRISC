`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Nick Markels
// 
// Create Date: 02/09/2023 03:46:21 PM
// Design Name: 
// Module Name: Data_path
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Data_path();


//Parameters
parameter DWIDTH = 32;

wire rd_addA, rd_addrB, wr_addr, wr_data;




endmodule
